LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY DFF8 IS 
	PORT(CLK: IN STD_LOGIC;
			WR:IN STD_LOGIC;
			D: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			Q: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END;
ARCHITECTURE ONE OF DFF8 IS
	SIGNAL S : STD_LOGIC_VECTOR(7 DOWNTO 0);
	BEGIN
		PROCESS (CLK,D,WR)
			BEGIN
				IF CLK'EVENT AND CLK = '1' THEN 
					IF WR = '1' THEN 
						S(7 DOWNTO 0) <= D(7 DOWNTO 0);
					END IF;
				END IF;
		END PROCESS;
Q(7 DOWNTO 0) <= S(7 DOWNTO 0);
END ONE;